Rsa256/synthesis/submodules/Rsa256Core.sv