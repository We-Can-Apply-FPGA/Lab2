Rsa256/synthesis/submodules/Rsa256Wrapper.sv